`timescale 1ns / 1ps

module CLA (
  input  logic [7:0] a,
  input  logic [7:0] b,
  input  logic       c_in,
  output logic [7:0] sum,
  output logic       c_out
);

endmodule
