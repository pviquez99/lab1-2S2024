`timescale 1ns / 1ps

module display_7_segmentos(
    input  logic [15:0] sw_pi,
    input  logic        boton_izquierda_pi,
    input  logic        boton_derecha_pi,
    output logic [6:0]  LED_o
    );
    
endmodule
